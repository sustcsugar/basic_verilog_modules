module sp_sram
#(
    DEPTH = 1024,
    AWIDTH = 10,
    DWIDTH = 8,
)
(

);

endmodule


module dp_sram
#(
    DEPTH = 1024,
    AWIDTH = 10,
    DWIDTH = 8,
)
(

);

endmodule


module sp_sram
#(
    DEPTH = 1024,
    AWIDTH = 10,
    DWIDTH = 8,
)
(

);

endmodule

